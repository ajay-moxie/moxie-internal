** Profile: "SCHEMATIC1-bias"  [ C:\ORCAD\ORCAD_16.5_LITE\PROJECTS\Hi-Lo CutOut schematic\6v hilo cutout-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.5_Lite\tools\pspice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\SCHEMATIC1.net" 


.END
