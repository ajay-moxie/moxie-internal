** Profile: "SCHEMATIC1-DCanalysis"  [ D:\personal\LEDs\PROJECTS\leddriver-pspicefiles\schematic1\dcanalysis.sim ] 

** Creating circuit file "DCanalysis.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/personal/LEDs/models/osram/osram-5mmradial.lib" 
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.5_Lite\tools\pspice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10000ns 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
